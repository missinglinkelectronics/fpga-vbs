`resetall
`default_nettype none
`timescale 1 ns / 1 ps


module <FPGA_TOP> ();
endmodule


`resetall
